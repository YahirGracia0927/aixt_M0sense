// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fabián A. Rojas Acosta, Alberto Pinzón Valero and Fernando Martínez Santa
// Date: 2024
// License: MIT
//
// Description: UART module (Arduino Nano - ATmega328P port)
module uart

// #include "//wsl.localhost/Ubuntu-22.04/home/yago/M0sense_BL702_example/bl_mcu_sdk/drivers/bl702_driver/hal_drv/inc/hal_uart.h"
#include <hal_uart.h>